module hello_world;
	initial
		begin
			$display("hello gtkwave!");
			$finish;
		end
endmodule
